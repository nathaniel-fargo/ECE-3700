module Test1(
	input hey,
	output alsoHey
	);
	
	assign alsoHey = hey;
	
	
endmodule