module Top;

endmodule