module TestBench;

	reg [1:0] A;
	reg [1:0] B;
	reg [1:0] I;
	wire [1:0] F;
	
	reg [3:0] num;
	

	Structural1 struct_inst (
		.A(A),
		.B(B),
		.I(I),
		.F(F)
	);
	
	
	initial begin
	
		num = 4'h0;
	
		
		A = num[3:2];
		B = num[1:0];
	
		I = 2'b00;
		#5;
		I = 2'b01;
		#5;
		I = 2'b10;
		#5;
		I = 2'b11;
		#5;
		
		num = num + 1;
			
	end
endmodule